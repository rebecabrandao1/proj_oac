/*o que foi adicionado:
1 -  módulo hazardunit - identifica os riscos e gera os sinais de controle para evitá-los
2 -  sinais de controle adicionais na controller e datapath (PCSrcE) e também havia a existencia de sinais na riscv que não estavam sendo usados pois não havia o hazardunit (ResultSrcEb0, ForwardAE, ForwardBE, StallF, StallD, FlushD, FlushE, Rs1D, Rs2D, Rs1E, Rs2E, RdE, RdM, RdW, RegWriteM, RegWriteW)
*/
/* como funciona no datapath: O hazardunit é o componente central que observa as instruções, detecta dependências e gera os sinais de Forward (adiantar), Stall (pausar) e Flush (limpar) para garantir que o fluxo de execução no pipeline seja sempre correto.*/
/* O endereço que está no pc é usado para ler a instrução da memória no imem. A instrução vai ser lida e salva no pipeline do reg if/id. Essa instrução forne os números dos registradores relacionados, cujo o id vai decodificar. São lidos dos registradores: o imediato e o regfile. Esses valores lidos são armazenados no pipe de id/ex*/
/* Agora entra a parte do hazard detection: onde occoree o stall  avalia as instruções que estão sendo lidas no if/id e no id/ex. Se houver uma instrução de load na ex que está tentando usar um registrador que está sendo carregado, a unidade de hazard detecta isso e gera sinais de stall para pausar o pipeline. Isso impede que a próxima instrução avance até que os dados necessários estejam disponíveis, masntendo as instruções no mesmo lugar e força os campos de controle a estarem em 0.*/
/*Em suma,  se no mux de entrada da alu, o dado que vem do banco de registradores (regfile) for igual ao dado que está sendo carregado na memória (dmem), o hazardunit detecta isso e gera um stall para pausar o pipeline até que o dado esteja disponível. Isso evita que a alu use um valor incorreto ou desatualizado, garantindo a integridade dos dados e a correta execução das instruções no pipeline.*/
/*Sobre a execuçaõ e o forwarding: é onde a alu opera (agora a instrução armazenada no id/ex é enviada para a lu que possui dois multiplexadores de entrada controlados pela unidade de fowarding que detecta se o operando que a alu precisa está disponível e m um operador de pipeline (ex/mem mem/wb) e ainda não foi escrito de volta no regfile. Se estiver disponível, o mux seleciona esse valor para a alu, caso contrário, seleciona o valor do regfile. Isso permite que a alu use os dados mais recentes sem esperar que sejam escritos de volta no regfile, melhorando a eficiência do pipeline e reduzindo stalls desnecessários.*/)
/* Os sinais forward a e forward b são usados para direcionar os multiplexadores que escolhem os dados para alu (como o valor encaminhado de ex/mem ou mem/wb). A alu vai executar o cálculo para load/store*/
/* Na fase de memória o resultado da alu é colcoado no reg ex/mem, se a instrução for um store, os dados a serem escritos na memória são provenientes do regfile (que podem ter sido encaminhados se necessário). Se for um load, os dados lidos da memória são armazenados no pipeline mem/wb.*/
/* Por fim, a escrita de volta WB os dados da alu ou os lidos da memória são escritos de volta no regfile e lido em MEM/WB  garantindo que o número de registrador de destino coreeto é passado e que seja usado, completando o ciclo de execução da instrução.*/
module hazardunit(input  logic        clk, reset,
                    input  logic [4:0]  Rs1D, Rs2D, Rs1E, Rs2E, RdE, RdM, RdW,
                    input  logic        RegWriteM, RegWriteW,
                    input  logic        ResultSrcEb0,
                    input  logic        PCSrcE,        // ADICIONADO: sinal de controle de desvio/jump
                    output logic [1:0]  ForwardAE, ForwardBE,
                    output logic        StallF, StallD, FlushD, FlushE);

/*entradas: clk, reset, Rs1D, Rs2D, Rs1E, Rs2E, RdE, RdM, RdW, RegWriteM, RegWriteW, ResultSrcEb0
saídas: ForwardAE, ForwardBE, StallF, StallD, FlushD, FlushE
Rs1D, Rs2D: registradores de origem na fase de decodificação (ID)
Rs1E, Rs2E: registradores de origem na fase de execução (EX)  */
/* o always_comb abaixo implementa a lógica para o encadeamento (forwarding) dos dados para a entrada A da ALU (ForwardAE).
Se a instrução na fase de memória (MEM) está escrevendo em um registrador (RegWriteM) e o registrador de destino (RdM) é igual ao registrador de origem 1 na fase de execução (Rs1E), então os dados são encaminhados da fase MEM (ForwardAE = 2'b10).
Se a instrução na fase de escrita (WB) está escrevendo em um registrador (RegWriteW) e o registrador de destino (RdW) é igual ao registrador de origem 1 na fase de execução (Rs1E), então os dados são encaminhados da fase WB (ForwardAE = 2'b01).
Caso contrário, os dados são usados diretamente da fase de decodificação (ForwardAE = 2'b00).*/
  always_comb
    if (RegWriteM & (RdM != 0) & (RdM == Rs1E))
      ForwardAE = 2'b10; // from MEM stage  -- o primeiro comando da Alu vem encaminhado de alguma operação anterior da alu
    else if (RegWriteW & (RdW != 0) & (RdW == Rs1E))
      ForwardAE = 2'b01; // from WB stage -- o primeiro comando da Alu vem encaminhado da memória de dados ou de alguma operação anterior da alu
    else
      ForwardAE = 2'b00; // from ID/EX stage -- o primeiro comando da Alu vem do banco de registradores

  // similar ao anterior, mas para a entrada B da ALU (ForwardBE)
  always_comb
    if (RegWriteM & (RdM != 0) & (RdM == Rs2E))
      ForwardBE = 2'b10; // from MEM stage  -- o segundo comando da Alu vem encaminhado de alguma operação anterior da alu
    else if (RegWriteW & (RdW != 0) & (RdW == Rs2E))
      ForwardBE = 2'b01; // from WB stage -- o segundo operando da Alu vem encaminhado da memória de dados ou de alguma operação anterior da alu
    else
      ForwardBE = 2'b00; // from ID/EX stage o segundo operando da Alu vem do banco de registradores
/*Além disso, o hazardunit também detecta as situações que envolve stalls e flushes:
- StallF e StallD são ativados quando há um risco de dados devido a uma instrução de carregamento (load) na fase de execução (EX) que está tentando usar um registrador que está sendo carregado. Isso é indicado por ResultSrcEb0 (que indica que a instrução atual na fase EX é um load) e a comparação dos registradores Rs1D e Rs2D com RdE.
- FlushD é ativado quando há um desvio (branch) ou salto (jump) na fase de execução (EX), indicado por PCSrcE.
- FlushE é ativado tanto por stalls (StallF) quanto por desvios/jumps (PCSrcE). Isso garante que a instrução na fase de execução seja descartada se houver um desvio ou se houver um stall necessário.    
*/

  assign StallF = (ResultSrcEb0 & ((RdE == Rs1D) | (RdE == Rs2D))) ? 1 : 0; // se a instrução na fase EX é um load e o registrador de destino (RdE) é igual a qualquer um dos registradores de origem na fase ID (Rs1D ou Rs2D), então StallF é ativado
  assign StallD = StallF; // StallD é ativado nas mesmas condições que StallF
  assign FlushD = PCSrcE; // FlushD é ativado se houver um desvio ou salto na fase EX
  assign FlushE = StallF || PCSrcE; // PCSrcE needs to be defined in the context where hazardunit is used
endmodule

module top(input  logic        clk, reset,  /*module top(): funciona como uma main, faz as chamadas dos demais módulos e integra CPU single-cycle RISC-V, memória de instruções e memória de dados [imem() e dmem()] e o hazardunit. entradas: clk, reset, WriteDataM; saídas: WriteDataM, DataAdrM, MemWriteM */
           output logic [31:0] WriteDataM, DataAdrM,  
           output logic        MemWriteM);

  logic [31:0] PCF, InstrF, ReadDataM; /* sinais de controle para o hazard unit */
  
  // instantiate processor and memories
  riscv riscv(clk, reset, PCF, InstrF, MemWriteM, DataAdrM,  /*instanciando o processador riscv, passando os sinais de controle e os sinais de entrada/saída*/
              WriteDataM, ReadDataM);
  imem imem(PCF, InstrF); /*instanciando a memória de instruções, passando o endereço do programa (PCF) e recebendo a instrução (InstrF)*/
  dmem dmem(clk, MemWriteM, DataAdrM, WriteDataM, ReadDataM); /*instanciando a memória de dados, passando o sinal de controle de escrita (MemWriteM), o endereço dos dados (DataAdrM), os dados a serem escritos (WriteDataM) e recebendo os dados lidos (ReadDataM)*/
endmodule

module riscv(input  logic        clk, reset,  /*module riscv(): implementa uma CPU RISC-V de 5 estágios com pipeline. entradas: clk, reset; saídas: PCF, InstrF, MemWriteM, ALUResultM, WriteDataM; entradas: ReadDataM */
             output logic [31:0] PCF,
             input  logic [31:0] InstrF,
             output logic        MemWriteM,
             output logic [31:0] ALUResultM, WriteDataM,
             input  logic [31:0] ReadDataM);

  logic [6:0]  opD;
  logic [2:0]  funct3D;
  logic        funct7b5D;
  logic [1:0]  ImmSrcD;
  logic        ZeroE;
  logic        PCSrcE;
  logic [2:0]  ALUControlE;
  logic        ALUSrcE;
  logic 	   ResultSrcEb0;
  logic        RegWriteM;
  logic [1:0]  ResultSrcW;
  logic        RegWriteW;

  logic [1:0]  ForwardAE, ForwardBE;
  logic        StallF, StallD, FlushD, FlushE;

  logic [4:0] Rs1D, Rs2D, Rs1E, Rs2E, RdE, RdM, RdW;

  controller c(clk, reset,  /*o controller chama os sinais de datapath, hazardunit e controller*/
               opD, funct3D, funct7b5D, ImmSrcD,
               FlushE, ZeroE, PCSrcE, ALUControlE, ALUSrcE, ResultSrcEb0,
               MemWriteM, RegWriteM, 
			   RegWriteW, ResultSrcW);

  hazardunit hu(clk, reset,
                Rs1D, Rs2D, Rs1E, Rs2E, RdE, RdM, RdW,
                RegWriteM, RegWriteW, ResultSrcEb0, PCSrcE,
                ForwardAE, ForwardBE, StallF, StallD, FlushD, FlushE);

  datapath dp(clk, reset,
              StallF, PCF, InstrF,
			  opD, funct3D, funct7b5D, StallD, FlushD, ImmSrcD,
			  FlushE, ForwardAE, ForwardBE, PCSrcE, ALUControlE, ALUSrcE, ZeroE,
              MemWriteM, WriteDataM, ALUResultM, ReadDataM,
              RegWriteW, ResultSrcW,
              Rs1D, Rs2D, Rs1E, Rs2E, RdE, RdM, RdW);

endmodule


module controller(input  logic		 clk, reset, // o módulo controller gera os sinais de controle necessários para o funcionamento do processador RISC-V, coordenando as operações em diferentes estágios do pipeline.
                  // Decode stage control signals  //entradas: opD(opcode) que pega os últimos 6 bits de Instr. funct3D: complemento de 3 bits do opcode, funct7b5: É o bit 5 do function7 (complemento de 7 bits do opcode), FlushE, Zero: Flag que vem da ALU e determina se branch de beq deve ser atendido. se  =1 o branch é atendido. Os sinais com D no final são da fase de decodificação, com E são da fase de execução, com M são da fase de memória e com W são da fase de escrita.
                  input logic [6:0]  opD,
                  input logic [2:0]  funct3D,
                  input logic 	     funct7b5D,
                  output logic [1:0] ImmSrcD,
                  // Execute stage control signals
                  input logic 	     FlushE, 
                  input logic 	     ZeroE, 
                  output logic       PCSrcE,        // for datapath and Hazard Unit
                  output logic [2:0] ALUControlE, 
                  output logic 	     ALUSrcE,
                  output logic       ResultSrcEb0,  // for Hazard Unit
                  // Memory stage control signals
                  output logic 	     MemWriteM,
                  output logic       RegWriteM,     // for Hazard Unit				  
                  // Writeback stage control signals
                  output logic 	     RegWriteW,     // for datapath and Hazard Unit
                  output logic [1:0] ResultSrcW);

  // pipelined control signals
  logic 	  RegWriteD, RegWriteE;
  logic [1:0] ResultSrcD, ResultSrcE, ResultSrcM;
  logic       MemWriteD, MemWriteE;
  logic		  JumpD, JumpE;
  logic		  BranchD, BranchE;
  logic	[1:0] ALUOpD;
  logic [2:0] ALUControlD;
  logic 	  ALUSrcD;
	
  // Decode stage logic
  maindec md(opD, ResultSrcD, MemWriteD, BranchD,
             ALUSrcD, RegWriteD, JumpD, ImmSrcD, ALUOpD);
  aludec  ad(opD[5], funct3D, funct7b5D, ALUOpD, ALUControlD);
  
  // Execute stage pipeline control register and logic
  floprc #(10) controlregE(clk, reset, FlushE,
                           {RegWriteD, ResultSrcD, MemWriteD, JumpD, BranchD, ALUControlD, ALUSrcD},
                           {RegWriteE, ResultSrcE, MemWriteE, JumpE, BranchE, ALUControlE, ALUSrcE});

  assign PCSrcE = (BranchE & ZeroE) | JumpE;
  assign ResultSrcEb0 = ResultSrcE[0];
  
  // Memory stage pipeline control register
  flopr #(4) controlregM(clk, reset,
                         {RegWriteE, ResultSrcE, MemWriteE},
                         {RegWriteM, ResultSrcM, MemWriteM});
  
  // Writeback stage pipeline control register
  flopr #(3) controlregW(clk, reset,
                         {RegWriteM, ResultSrcM},
                         {RegWriteW, ResultSrcW});     
endmodule

module maindec(input  logic [6:0] op,
               output logic [1:0] ResultSrc,
               output logic       MemWrite,
               output logic       Branch, ALUSrc,
               output logic       RegWrite, Jump,
               output logic [1:0] ImmSrc,
               output logic [1:0] ALUOp);

  logic [10:0] controls;

  assign {RegWrite, ImmSrc, ALUSrc, MemWrite,
          ResultSrc, Branch, ALUOp, Jump} = controls;

  always_comb
    case(op)
    // RegWrite_ImmSrc_ALUSrc_MemWrite_ResultSrc_Branch_ALUOp_Jump
      7'b0000011: controls = 11'b1_00_1_0_01_0_00_0; // lw
      7'b0100011: controls = 11'b0_01_1_1_00_0_00_0; // sw
      7'b0110011: controls = 11'b1_xx_0_0_00_0_10_0; // R-type 
      7'b1100011: controls = 11'b0_10_0_0_00_1_01_0; // beq
      7'b0010011: controls = 11'b1_00_1_0_00_0_10_0; // I-type ALU
      7'b1101111: controls = 11'b1_11_0_0_10_0_00_1; // jal
      7'b0000000: controls = 11'b0_00_0_0_00_0_00_0; // need valid values at reset
      default:    controls = 11'bx_xx_x_x_xx_x_xx_x; // non-implemented instruction
    endcase
endmodule

module aludec(input  logic       opb5,
              input  logic [2:0] funct3,
              input  logic       funct7b5, 
              input  logic [1:0] ALUOp,
              output logic [2:0] ALUControl);

  logic  RtypeSub;
  assign RtypeSub = funct7b5 & opb5;  // TRUE for R-type subtract instruction

  always_comb
    case(ALUOp)
      2'b00:                ALUControl = 3'b000; // addition
      2'b01:                ALUControl = 3'b001; // subtraction
      default: case(funct3) // R-type or I-type ALU
                 3'b000:  if (RtypeSub) 
                            ALUControl = 3'b001; // sub
                          else          
                            ALUControl = 3'b000; // add, addi
                 3'b010:    ALUControl = 3'b101; // slt, slti
                 3'b110:    ALUControl = 3'b011; // or, ori
                 3'b111:    ALUControl = 3'b010; // and, andi
                 default:   ALUControl = 3'bxxx; // ???
               endcase
    endcase
endmodule

module datapath(input logic clk, reset,
                // Fetch stage signals
                input  logic        StallF,
                output logic [31:0] PCF,
                input  logic [31:0] InstrF,
                // Decode stage signals
                output logic [6:0]  opD,
                output logic [2:0]	funct3D, 
                output logic        funct7b5D,
                input  logic        StallD, FlushD,
                input  logic [1:0]  ImmSrcD,
                // Execute stage signals
                input  logic        FlushE,
                input  logic [1:0]  ForwardAE, ForwardBE,
                input  logic        PCSrcE,
                input  logic [2:0]  ALUControlE,
                input  logic        ALUSrcE,
                output logic        ZeroE,
                // Memory stage signals
                input  logic        MemWriteM, 
                output logic [31:0] WriteDataM, ALUResultM,
                input  logic [31:0] ReadDataM,
                // Writeback stage signals
                input  logic        RegWriteW, 
                input  logic [1:0]  ResultSrcW,
                // Hazard Unit signals 
                output logic [4:0]  Rs1D, Rs2D, Rs1E, Rs2E,
                output logic [4:0]  RdE, RdM, RdW);

  // Fetch stage signals
  logic [31:0] PCNextF, PCPlus4F;
  // Decode stage signals
  logic [31:0] InstrD;
  logic [31:0] PCD, PCPlus4D;
  logic [31:0] RD1D, RD2D;
  logic [31:0] ImmExtD;
  logic [4:0]  RdD;
  // Execute stage signals
  logic [31:0] RD1E, RD2E;
  logic [31:0] PCE, ImmExtE;
  logic [31:0] SrcAE, SrcBE;
  logic [31:0] ALUResultE;
  logic [31:0] WriteDataE;
  logic [31:0] PCPlus4E;
  logic [31:0] PCTargetE;
  // Memory stage signals
  logic [31:0] PCPlus4M;
  // Writeback stage signals
  logic [31:0] ALUResultW;
  logic [31:0] ReadDataW;
  logic [31:0] PCPlus4W;
  logic [31:0] ResultW;

  // Fetch stage pipeline register and logic
  mux2    #(32) pcmux(PCPlus4F, PCTargetE, PCSrcE, PCNextF);
  flopenr #(32) pcreg(clk, reset, ~StallF, PCNextF, PCF);
  adder         pcadd(PCF, 32'h4, PCPlus4F);

  // Decode stage pipeline register and logic
  flopenrc #(96) regD(clk, reset, FlushD, ~StallD, 
                      {InstrF, PCF, PCPlus4F},
                      {InstrD, PCD, PCPlus4D});
  assign opD       = InstrD[6:0];
  assign funct3D   = InstrD[14:12];
  assign funct7b5D = InstrD[30];
  assign Rs1D      = InstrD[19:15];
  assign Rs2D      = InstrD[24:20];
  assign RdD       = InstrD[11:7];
	
  regfile        rf(clk, RegWriteW, Rs1D, Rs2D, RdW, ResultW, RD1D, RD2D);
  extend         ext(InstrD[31:7], ImmSrcD, ImmExtD);
 
  // Execute stage pipeline register and logic
  floprc #(175) regE(clk, reset, FlushE, 
                     {RD1D, RD2D, PCD, Rs1D, Rs2D, RdD, ImmExtD, PCPlus4D}, 
                     {RD1E, RD2E, PCE, Rs1E, Rs2E, RdE, ImmExtE, PCPlus4E});
	
  mux3   #(32)  faemux(RD1E, ResultW, ALUResultM, ForwardAE, SrcAE);
  mux3   #(32)  fbemux(RD2E, ResultW, ALUResultM, ForwardBE, WriteDataE);
  mux2   #(32)  srcbmux(WriteDataE, ImmExtE, ALUSrcE, SrcBE);
  alu           alu(SrcAE, SrcBE, ALUControlE, ALUResultE, ZeroE);
  adder         branchadd(ImmExtE, PCE, PCTargetE);

  // Memory stage pipeline register
  flopr  #(101) regM(clk, reset, 
                     {ALUResultE, WriteDataE, RdE, PCPlus4E},
                     {ALUResultM, WriteDataM, RdM, PCPlus4M});
	
  // Writeback stage pipeline register and logic
  flopr  #(101) regW(clk, reset, 
                     {ALUResultM, ReadDataM, RdM, PCPlus4M},
                     {ALUResultW, ReadDataW, RdW, PCPlus4W});
  mux3   #(32)  resultmux(ALUResultW, ReadDataW, PCPlus4W, ResultSrcW, ResultW);	
endmodule


module regfile(input  logic        clk, 
               input  logic        we3, 
               input  logic [ 4:0] a1, a2, a3, 
               input  logic [31:0] wd3, 
               output logic [31:0] rd1, rd2);

  logic [31:0] rf[31:0];

  // three ported register file
  // read two ports combinationally (A1/RD1, A2/RD2)
  // write third port on rising edge of clock (A3/WD3/WE3)
  // write occurs on falling edge of clock
  // register 0 hardwired to 0

  always_ff @(negedge clk)
    if (we3) rf[a3] <= wd3;	

  assign rd1 = (a1 != 0) ? rf[a1] : 0;
  assign rd2 = (a2 != 0) ? rf[a2] : 0;
endmodule

module adder(input  [31:0] a, b,
             output [31:0] y);

  assign y = a + b;
endmodule

module extend(input  logic [31:7] instr,
              input  logic [1:0]  immsrc,
              output logic [31:0] immext);
 
  always_comb
    case(immsrc) 
               // I-type 
      2'b00:   immext = {{20{instr[31]}}, instr[31:20]};  
               // S-type (stores)
      2'b01:   immext = {{20{instr[31]}}, instr[31:25], instr[11:7]}; 
               // B-type (branches)
      2'b10:   immext = {{20{instr[31]}}, instr[7], instr[30:25], instr[11:8], 1'b0}; 
               // J-type (jal)
      2'b11:   immext = {{12{instr[31]}}, instr[19:12], instr[20], instr[30:21], 1'b0}; 
      default: immext = 32'bx; // undefined
    endcase             
endmodule

module flopr #(parameter WIDTH = 8) // o módulo flopr é um flip-flop com reset assíncrono
              (input  logic             clk, reset, //entradas: clk: clock, reset: controle do flip flop, d: informação do estado final
               input  logic [WIDTH-1:0] d,  
               output logic [WIDTH-1:0] q); //saídas: q: informação do estado inicial

  always_ff @(posedge clk, posedge reset) ///mudanças de estados só acontecem baseadas no clik e reset
    if (reset) q <= 0; //se reset=1, é necessario apagar a informação do flipflop, entao a saida é 0 e não armazena nada no pc
    else       q <= d; //// caso contrário, q recebe a informação do estadoa tual
endmodule

module flopenr #(parameter WIDTH = 8)
                (input  logic             clk, reset, en,
                 input  logic [WIDTH-1:0] d, 
                 output logic [WIDTH-1:0] q);

  always_ff @(posedge clk, posedge reset)
    if (reset)   q <= 0;
    else if (en) q <= d;
endmodule

module flopenrc #(parameter WIDTH = 8) // o módulo flopenrc é um flip-flop com sinal de habilitação e limpeza assíncrona
                (input  logic             clk, reset, clear, en, //entradas: clk: clock, reset: sinal de reset assíncrono, clear: sinal de limpeza assíncrona, en: sinal de habilitação, d: dado de entrada de WIDTH bits
                 input  logic [WIDTH-1:0] d, 
                 output logic [WIDTH-1:0] q); //saídas: q: dado de saída de WIDTH bits

  always_ff @(posedge clk, posedge reset) //ação que sempre acontecerá na saída do clock ou no reset
    if (reset)   q <= 0; //se reset for igual a 1 , q recebe 0
    else if (en)  //se en for igual a 1 , q recebe o valor de d
      if (clear) q <= 0; //se clear for igual a 1 , q recebe 0
      else       q <= d; //se clear for igual a 0 , q recebe o valor de d
endmodule

module floprc #(parameter WIDTH = 8) // o módulo floprc é um flip-flop com sinal de limpeza assíncrona
              (input  logic clk, //entradas: clk: clock, reset: sinal de reset assíncrono, clear: sinal de limpeza assíncrona, d: dado de entrada de WIDTH bits
               input  logic reset,
               input  logic clear,
               input  logic [WIDTH-1:0] d, 
               output logic [WIDTH-1:0] q); //saídas: q: dado de saída de WIDTH bits

  always_ff @(posedge clk, posedge reset) //ação que sempre acontecerá na saída do clock ou no reset
    if (reset) q <= 0; //se reset for igual a 1 , q recebe 0
    else       
      if (clear) q <= 0; //se clear for igual a 1 , q recebe 0
      else       q <= d; //se clear for igual a 0 , q recebe o valor de d
endmodule

module mux2 #(parameter WIDTH = 8) // multiplexador de 2 entradas
             (input  logic [WIDTH-1:0] d0, d1, // entradas: d0, d1: dados de entrada de WIDTH bits
              input  logic             s, // seletor para escolher entre as 2 entradas
              output logic [WIDTH-1:0] y); // saídas: y: dado de saída de WIDTH bits

  assign y = s ? d1 : d0; 
endmodule

module mux3 #(parameter WIDTH = 8) // multiplexador de 3 entradas
             (input  logic [WIDTH-1:0] d0, d1, d2, // entradas: d0, d1, d2: dados de entrada de WIDTH bits
              input  logic [1:0]       s, // seletor de 2 bits para escolher entre as 3 entradas
              output logic [WIDTH-1:0] y); // saídas: y: dado de saída de WIDTH bits

  assign y = s[1] ? d2 : (s[0] ? d1 : d0); // se s[1] for 1, y recebe d2; se s[1] for 0 e s[0] for 1, y recebe d1; caso contrário, y recebe d0 
endmodule

module imem(input  logic [31:0] a,  //entradas: a instrução de 32 bits que representa o PC
            output logic [31:0] rd); //saídas: rd devolve a instrução lida

  logic [31:0] RAM[63:0]; //memória do computador (uma matriz 64 linhas de 32 bits)

  initial
      $readmemh("riscvtest.txt",RAM); //lê o arquivo de teste

  assign rd = RAM[a[31:2]]; // word aligned // word aligned recebe todas as linhas com os bits de 2 a 31
endmodule

module dmem(input  logic        clk, we,  //entradas clock, we:sinal para fazer a escrita da informação recebida por a , a:saida obtida pela ULA que pode variar de endereços a resultado de contas, wd:dado recebido pelo Register File (regfile),
            input  logic [31:0] a, wd,
            output logic [31:0] rd); //saídas: rd:ReadData: Quando a=endereço de memória rd é o dado que esse endereço carrega logic [31:0] RAM[63:0]

  logic [31:0] RAM[63:0];

  assign rd = RAM[a[31:2]]; // word aligned

  always_ff @(posedge clk) //ação que sempre acontecerá na saída do clock
    if (we) RAM[a[31:2]] <= wd; //se MemoryWrite for igual a  1 , a inforação recebida na entrada "a" (vindo da ula) é escrita 
endmodule

module alu(input  logic [31:0] a, b,/*entradas: a, b: um valor a ser operado, alucontrol: um controle de 3 bits que vai definir a operação entre a e b; saídas:  //saídas: result: vai ser o resultadod de f(a,b), zero: Comparação entre a e b: se a=b, zero = 1 se nãp zero=0, condinvb: avalia se necessita inverter b para alguma operação, sum:resultado da soma v:verifica se tem overflow na operaçao, isaddSub: verifica qual operação é necessária se soma ou subtração*/
           input  logic [2:0]  alucontrol,
           output logic [31:0] result,
           output logic        zero);

  logic [31:0] condinvb, sum;
  logic        v;              // overflow
  logic        isAddSub;       // true when is add or subtract operation

  assign condinvb = alucontrol[0] ? ~b : b; //inverte os bits de b de acordo com o aluontrol se alucontrol[0]=1 a inversão é feita, caso contrário não.
  assign sum = a + condinvb + alucontrol[0];
  assign isAddSub = ~alucontrol[2] & ~alucontrol[1] |
                    ~alucontrol[1] &  alucontrol[0];

  always_comb
    case (alucontrol)
      3'b000:  result = sum;         // add
      3'b001:  result = sum;         // subtract
      3'b010:  result = a & b;       // and
      3'b011:  result = a | b;       // or
      3'b100:  result = a ^ b;       // xor
      3'b101:  result = sum[31] ^ v; // slt
      3'b110:  result = a << b[4:0]; // sll
      3'b111:  result = a >> b[4:0]; // srl
      default: result = 32'bx;
    endcase

  assign zero = (result == 32'b0);
  assign v = ~(alucontrol[0] ^ a[31] ^ b[31]) & (a[31] ^ sum[31]) & isAddSub;
  
endmodule